/*
forwarding unit module
*/

// interface include
`include "forwarding_unit_if.vh"
// memory types
`include "cpu_types_pkg.vh"

module forwarding_unit (
  forwarding_unit_if.fu fuif
);




always_comb begin

end

endmodule
